// SPI Interface
interface spi_if(input logic clk, rst);
    logic mosi, miso, sck, ss;
endinterface