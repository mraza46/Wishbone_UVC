package my_package;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "wb_seq_item.sv"
  `include "wb_seq.sv"
  `include "wb_sequencer.sv"
  `include "wb_driver.sv"
  `include "wb_monitor.sv"
  `include "wb_agent.sv"
  //`include "wb_scoreboard.sv"
  `include "wb_env.sv"
  `include "wb_test.sv"

endpackage

